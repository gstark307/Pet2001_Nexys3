`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////
//
// Engineer:         Thomas Skibo
// 
// Create Date:      Aug 24, 2011
//
// Module Name:      Pet2001_Nexys3
//
// Target Devices:   Xilinx Spartan-6 XC6SLX16
//
// Description:     Top module for Commodore Pet emulator on Digilent Nexys3
//                  Spartan 6 evaluation board.  I/O's at this level represent
//		    pins on the Spartan 6.
//
// Additional Comments:
//
//	Nexys3 I/O assigns:
//
//		SW[0] -	Full speed CPU clocking (vs. 100-to-1 slowdown)
//		SW[1] -	Stop CPU
//		SW[2] -	Diag (connected to PORTA[7] of PIA1)
//		SW[3] - Cassette Sense
//
//		btns -	Full reset
//
//		Led[0] - Cassette Write
//		Led[1] - Cassette Motor
//		Led[2] - Audio
//		Led[3] - RS232 CTS#
//
//		JA[3] -	RS232 CTS# (output: need to wire to FT232)
//		JA[4] -	Keyboard PS2 Clock (input)
//		JA[6] -	Keyboard PS2 Data (input)
//
//		JB[0] -	Audio
//		JB[1] -	Cassette Data Write (output)
//		JB[2] -	Cassette Data Read (output - generated by cass232)
//		JB[3] - Cassette Motor
//
//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2011, Thomas Skibo.  All rights reserved.
// 
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
// * Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.
// * Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.
// * The names of contributors may not be used to endorse or promote products
//   derived from this software without specific prior written permission.
// 
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL Thomas Skibo OR CONTRIBUTORS BE LIABLE FOR
// ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE
// USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
//////////////////////////////////////////////////////////////////////////////

module pet2001(	input          		btns,		// Buttons
		input			btnu,
		input			btnl,
		input			btnd,
		input			btnr,

		input  [7:0]   		sw,		// Switches

		output reg [7:0]	Led,		// LEDs

		output [2:0]   		vgaRed,
		output [2:0]   		vgaGreen,
		output [2:1]   		vgaBlue,
		output         		Hsync,
		output         		Vsync,

		input			Rs232RxD,
		output			Rs232TxD,

		output [7:0]   		seg,		// 7-seg disp cathodes
		output [3:0]   		an,		// 7-seg disp anodes

		inout [7:0]		JA,		// 12-pin PMOD conn
		inout [7:0]		JB,		// 12-pin PMOD conn

		input          		clk_100M	// 100 Mhz clock
	);

`ifdef simulation
 `include "roms/pet2001_rom1.v"
`endif

   //////////////////////////////////////////////////////////////////////
   // Create global clock and synchronous system reset.                //
   //////////////////////////////////////////////////////////////////////

    wire 	clknub;
    wire 	clk;
    wire 	locked;

    // Use DCM.
    DCM_SP #(.CLKIN_PERIOD(10.000),
	     .CLKIN_DIVIDE_BY_2("true"))
    	DCM_SP_INST (
                     .CLKIN(clk_100M),
                     .CLKFB(clk),
                     .RST(1'b0),
                     .PSEN(1'b0),
                     .PSINCDEC(1'b0),
                     .PSCLK(1'b0),
                     .DSSEN(1'b0),
                     .CLK0(clknub),
                     .CLK90(),
                     .CLK180(),
                     .CLK270(),
                     .CLKDV(),
                     .CLK2X(),
                     .CLK2X180(),
                     .CLKFX(),
                     .CLKFX180(),
                     .STATUS(),
                     .LOCKED(locked),
                     .PSDONE()
	     );

    // Put clk on clock network.
    BUFG BG (.I(clknub), .O(clk));

    // Synchronize reset.
    wire 	reset_unsynced = ! locked || btns;
    wire 	reset_unsynced_1;
    wire 	reset;
   
    FDP #(.INIT(1'b1)) sync_reset_1(.Q(reset_unsynced_1),
				    .D(reset_unsynced),
				    .C(clk),
				    .PRE(1'b0));
    FDP #(.INIT(1'b1)) sync_reset_2(.Q(reset),
				    .D(reset_unsynced_1),
				    .C(clk),
				    .PRE(1'b0));

    ////////////////////////////////////////////////////////////////////////
    // Synchronize switch inputs
    ////////////////////////////////////////////////////////////////////////
    reg [7:0] 	sw_1;
    reg [7:0] 	sw_2;
    always @(posedge clk)
	if (reset) begin
            sw_1 <= 8'd0;
            sw_2 <= 8'd0;
	end
	else begin
            sw_1 <= sw;
            sw_2 <= sw_1;
	end

    wire diag_l = ~sw_2[2];
    wire clk_stop = sw_2[1];
    wire clk_speed = sw_2[0];

    /////////////////////////////////////////////////////////////////////
    // Top level module
    /////////////////////////////////////////////////////////////////////

    wire [2:0]	vgaBlueAll;
    assign	vgaBlue = vgaBlueAll[2:1];
    
    wire 	ps2_clk = JA[4];
    wire 	ps2_data = JA[6];
    
    wire [7:0] 	keyin;				// PET keyboard matrix
    wire [3:0] 	keyrow;
    
    wire 	cass_motor_n;
    wire 	cass_write;
    wire 	cass_sense_n = ~sw_2[3];
    wire 	cass_read;
    
    wire 	audio;

    pet2001_top pet_top(.vgaRed(vgaRed),
			.vgaGreen(vgaGreen),
			.vgaBlue(vgaBlueAll),
			.Hsync(Hsync),
			.Vsync(Vsync),

			.keyrow(keyrow),
			.keyin(keyin),
	
			.cass_motor_n(cass_motor_n),
			.cass_write(cass_write),
			.cass_sense_n(cass_sense_n),
			.cass_read(cass_read),
        
			.audio(audio),

			.diag_l(diag_l),
        
			.clk_speed(clk_speed),
			.clk_stop(clk_stop),

			.clk(clk),
			.reset(reset)
		);

    assign	JB[0] = audio;
    assign	JB[1] =	cass_write;
    assign	JB[2] =	cass_read;
    assign	JB[3] = ~cass_motor_n;

    //////////////////////////////////////////////////////////////////////
    // RS-232 to Cassette Interface
    //////////////////////////////////////////////////////////////////////

    wire        Rs232CtsN;
   
    pet2001cass232 cass(.tx232(Rs232TxD),
			.rx232(Rs232RxD),
			.cts232n(Rs232CtsN),

			.cass_motor_n(cass_motor_n),
			.cass_write(cass_write),
			.cass_read(cass_read),

			.clk(clk),
			.reset(reset)
		);

    assign JA[3] = Rs232CtsN;

    //////////////////////////////////////////////////////////////////////
    // PS/2 to PET keyboard interface
    //////////////////////////////////////////////////////////////////////

    pet2001ps2_key ps2key(.keyin(keyin),		// PET key matrix
			  .keyrow(keyrow),
			  
			  .ps2_clk(ps2_clk),		// PS/2 interface
			  .ps2_data(ps2_data),

			  .clk(clk),
			  .reset(reset)
		  );
	
    //////////////////////////////////////////////////////////////////////
    // Drive LEDs (could be more interesting).
    //////////////////////////////////////////////////////////////////////
    
    // Display mux
    dispmux dispmux0(.SevenSeg(seg),
                     .SevenAnode(an),

		     .dispA(8'b1010_0100),
		     .dispB(8'b1100_0000),
		     .dispC(8'b1100_0000),
		     .dispD(8'b1111_1001),

                     .reset(reset),
                     .clk(clk)
	     );

    always @(posedge clk)
	Led <= { 4'b0000, Rs232CtsN, audio, ~cass_motor_n, cass_write };
    
endmodule // pet2001

